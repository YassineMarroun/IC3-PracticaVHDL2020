--------------------------------
library IEEE;
use IEEE.std_logic_1164.all;

entity funcionF1F2 is
	port(F1, F2	:out std_logic;
	     x, y, z	:in std_logic);
end entity funcionF1F2;
--------------------------------